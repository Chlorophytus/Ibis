/**
 *  Copyright 2025 Roland Metivier
 *
 *  SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
 *
 *  Licensed under the Solderpad Hardware License v 2.1 (the "License"); you may
 *  not use this file except in compliance with the License, or, at your option,
 *  the Apache License version 2.0.
 *
 *  You may obtain a copy of the License at
 *
 *  https://solderpad.org/licenses/SHL-2.1/
 *
 *  Unless required by applicable law or agreed to in writing, any work
 *  distributed under the License is distributed on an "AS IS" BASIS, WITHOUT
 *  WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *
 *  See the License for the specific language governing permissions and
 *  limitations under the License.
 */
`timescale 1ns / 1ps
`default_nettype none
// AUTOGENERATED: 8-bit square root
module ibis_square_root
 (input wire logic unsigned [7:0] in_bits,
  output logic unsigned [7:0] square_root);
  always_comb begin: ibis_square_root_combinatorial
    unique case(in_bits) inside
      8'h00: square_root = 8'h00; // 0.0
      8'h01: square_root = 8'h10; // 1.0
      8'h02: square_root = 8'h16; // 1.4142135623730951
      8'h03: square_root = 8'h1B; // 1.7320508075688772
      8'h04: square_root = 8'h20; // 2.0
      8'h05: square_root = 8'h23; // 2.23606797749979
      8'h06: square_root = 8'h27; // 2.449489742783178
      8'h07: square_root = 8'h2A; // 2.6457513110645907
      8'h08: square_root = 8'h2D; // 2.8284271247461903
      8'h09: square_root = 8'h30; // 3.0
      8'h0A: square_root = 8'h32; // 3.1622776601683795
      8'h0B: square_root = 8'h35; // 3.3166247903554
      8'h0C: square_root = 8'h37; // 3.4641016151377544
      8'h0D: square_root = 8'h39; // 3.605551275463989
      8'h0E: square_root = 8'h3B; // 3.7416573867739413
      8'h0F: square_root = 8'h3D; // 3.872983346207417
      8'h10: square_root = 8'h40; // 4.0
      8'h11: square_root = 8'h41; // 4.123105625617661
      8'h12: square_root = 8'h43; // 4.242640687119285
      8'h13: square_root = 8'h45; // 4.358898943540674
      8'h14: square_root = 8'h47; // 4.47213595499958
      8'h15: square_root = 8'h49; // 4.58257569495584
      8'h16: square_root = 8'h4B; // 4.69041575982343
      8'h17: square_root = 8'h4C; // 4.795831523312719
      8'h18: square_root = 8'h4E; // 4.898979485566356
      8'h19: square_root = 8'h50; // 5.0
      8'h1A: square_root = 8'h51; // 5.0990195135927845
      8'h1B: square_root = 8'h53; // 5.196152422706632
      8'h1C: square_root = 8'h54; // 5.291502622129181
      8'h1D: square_root = 8'h56; // 5.385164807134504
      8'h1E: square_root = 8'h57; // 5.477225575051661
      8'h1F: square_root = 8'h59; // 5.5677643628300215
      8'h20: square_root = 8'h5A; // 5.656854249492381
      8'h21: square_root = 8'h5B; // 5.744562646538029
      8'h22: square_root = 8'h5D; // 5.830951894845301
      8'h23: square_root = 8'h5E; // 5.916079783099616
      8'h24: square_root = 8'h60; // 6.0
      8'h25: square_root = 8'h61; // 6.082762530298219
      8'h26: square_root = 8'h62; // 6.164414002968976
      8'h27: square_root = 8'h63; // 6.244997998398398
      8'h28: square_root = 8'h65; // 6.324555320336759
      8'h29: square_root = 8'h66; // 6.4031242374328485
      8'h2A: square_root = 8'h67; // 6.48074069840786
      8'h2B: square_root = 8'h68; // 6.557438524302
      8'h2C: square_root = 8'h6A; // 6.6332495807108
      8'h2D: square_root = 8'h6B; // 6.708203932499369
      8'h2E: square_root = 8'h6C; // 6.782329983125268
      8'h2F: square_root = 8'h6D; // 6.855654600401044
      8'h30: square_root = 8'h6E; // 6.928203230275509
      8'h31: square_root = 8'h70; // 7.0
      8'h32: square_root = 8'h71; // 7.0710678118654755
      8'h33: square_root = 8'h72; // 7.14142842854285
      8'h34: square_root = 8'h73; // 7.211102550927978
      8'h35: square_root = 8'h74; // 7.280109889280518
      8'h36: square_root = 8'h75; // 7.3484692283495345
      8'h37: square_root = 8'h76; // 7.416198487095663
      8'h38: square_root = 8'h77; // 7.483314773547883
      8'h39: square_root = 8'h78; // 7.54983443527075
      8'h3A: square_root = 8'h79; // 7.615773105863909
      8'h3B: square_root = 8'h7A; // 7.681145747868608
      8'h3C: square_root = 8'h7B; // 7.745966692414834
      8'h3D: square_root = 8'h7C; // 7.810249675906654
      8'h3E: square_root = 8'h7D; // 7.874007874011811
      8'h3F: square_root = 8'h7E; // 7.937253933193772
      8'h40: square_root = 8'h80; // 8.0
      8'h41: square_root = 8'h80; // 8.06225774829855
      8'h42: square_root = 8'h81; // 8.12403840463596
      8'h43: square_root = 8'h82; // 8.18535277187245
      8'h44: square_root = 8'h83; // 8.246211251235321
      8'h45: square_root = 8'h84; // 8.306623862918075
      8'h46: square_root = 8'h85; // 8.366600265340756
      8'h47: square_root = 8'h86; // 8.426149773176359
      8'h48: square_root = 8'h87; // 8.48528137423857
      8'h49: square_root = 8'h88; // 8.54400374531753
      8'h4A: square_root = 8'h89; // 8.602325267042627
      8'h4B: square_root = 8'h8A; // 8.660254037844387
      8'h4C: square_root = 8'h8B; // 8.717797887081348
      8'h4D: square_root = 8'h8C; // 8.774964387392123
      8'h4E: square_root = 8'h8D; // 8.831760866327848
      8'h4F: square_root = 8'h8E; // 8.888194417315589
      8'h50: square_root = 8'h8F; // 8.94427190999916
      8'h51: square_root = 8'h90; // 9.0
      8'h52: square_root = 8'h90; // 9.055385138137417
      8'h53: square_root = 8'h91; // 9.1104335791443
      8'h54: square_root = 8'h92; // 9.16515138991168
      8'h55: square_root = 8'h93; // 9.219544457292887
      8'h56: square_root = 8'h94; // 9.273618495495704
      8'h57: square_root = 8'h95; // 9.327379053088816
      8'h58: square_root = 8'h96; // 9.38083151964686
      8'h59: square_root = 8'h96; // 9.433981132056603
      8'h5A: square_root = 8'h97; // 9.486832980505138
      8'h5B: square_root = 8'h98; // 9.539392014169456
      8'h5C: square_root = 8'h99; // 9.591663046625438
      8'h5D: square_root = 8'h9A; // 9.643650760992955
      8'h5E: square_root = 8'h9B; // 9.695359714832659
      8'h5F: square_root = 8'h9B; // 9.746794344808963
      8'h60: square_root = 8'h9C; // 9.797958971132712
      8'h61: square_root = 8'h9D; // 9.848857801796104
      8'h62: square_root = 8'h9E; // 9.899494936611665
      8'h63: square_root = 8'h9F; // 9.9498743710662
      8'h64: square_root = 8'hA0; // 10.0
      8'h65: square_root = 8'hA0; // 10.04987562112089
      8'h66: square_root = 8'hA1; // 10.099504938362077
      8'h67: square_root = 8'hA2; // 10.14889156509222
      8'h68: square_root = 8'hA3; // 10.198039027185569
      8'h69: square_root = 8'hA3; // 10.246950765959598
      8'h6A: square_root = 8'hA4; // 10.295630140987
      8'h6B: square_root = 8'hA5; // 10.344080432788601
      8'h6C: square_root = 8'hA6; // 10.392304845413264
      8'h6D: square_root = 8'hA7; // 10.44030650891055
      8'h6E: square_root = 8'hA7; // 10.488088481701515
      8'h6F: square_root = 8'hA8; // 10.535653752852738
      8'h70: square_root = 8'hA9; // 10.583005244258363
      8'h71: square_root = 8'hAA; // 10.63014581273465
      8'h72: square_root = 8'hAA; // 10.677078252031311
      8'h73: square_root = 8'hAB; // 10.723805294763608
      8'h74: square_root = 8'hAC; // 10.770329614269007
      8'h75: square_root = 8'hAD; // 10.816653826391969
      8'h76: square_root = 8'hAD; // 10.862780491200215
      8'h77: square_root = 8'hAE; // 10.908712114635714
      8'h78: square_root = 8'hAF; // 10.954451150103322
      8'h79: square_root = 8'hB0; // 11.0
      8'h7A: square_root = 8'hB0; // 11.045361017187261
      8'h7B: square_root = 8'hB1; // 11.090536506409418
      8'h7C: square_root = 8'hB2; // 11.135528725660043
      8'h7D: square_root = 8'hB2; // 11.180339887498949
      8'h7E: square_root = 8'hB3; // 11.224972160321824
      8'h7F: square_root = 8'hB4; // 11.269427669584644
      8'h80: square_root = 8'hB5; // 11.313708498984761
      8'h81: square_root = 8'hB5; // 11.357816691600547
      8'h82: square_root = 8'hB6; // 11.40175425099138
      8'h83: square_root = 8'hB7; // 11.445523142259598
      8'h84: square_root = 8'hB7; // 11.489125293076057
      8'h85: square_root = 8'hB8; // 11.532562594670797
      8'h86: square_root = 8'hB9; // 11.575836902790225
      8'h87: square_root = 8'hB9; // 11.61895003862225
      8'h88: square_root = 8'hBA; // 11.661903789690601
      8'h89: square_root = 8'hBB; // 11.704699910719626
      8'h8A: square_root = 8'hBB; // 11.74734012447073
      8'h8B: square_root = 8'hBC; // 11.789826122551595
      8'h8C: square_root = 8'hBD; // 11.832159566199232
      8'h8D: square_root = 8'hBD; // 11.874342087037917
      8'h8E: square_root = 8'hBE; // 11.916375287812984
      8'h8F: square_root = 8'hBF; // 11.958260743101398
      8'h90: square_root = 8'hC0; // 12.0
      8'h91: square_root = 8'hC0; // 12.041594578792296
      8'h92: square_root = 8'hC1; // 12.083045973594572
      8'h93: square_root = 8'hC1; // 12.12435565298214
      8'h94: square_root = 8'hC2; // 12.165525060596439
      8'h95: square_root = 8'hC3; // 12.206555615733702
      8'h96: square_root = 8'hC3; // 12.24744871391589
      8'h97: square_root = 8'hC4; // 12.288205727444508
      8'h98: square_root = 8'hC5; // 12.328828005937952
      8'h99: square_root = 8'hC5; // 12.36931687685298
      8'h9A: square_root = 8'hC6; // 12.409673645990857
      8'h9B: square_root = 8'hC7; // 12.449899597988733
      8'h9C: square_root = 8'hC7; // 12.489995996796797
      8'h9D: square_root = 8'hC8; // 12.529964086141668
      8'h9E: square_root = 8'hC9; // 12.569805089976535
      8'h9F: square_root = 8'hC9; // 12.609520212918492
      8'hA0: square_root = 8'hCA; // 12.649110640673518
      8'hA1: square_root = 8'hCB; // 12.68857754044952
      8'hA2: square_root = 8'hCB; // 12.727922061357855
      8'hA3: square_root = 8'hCC; // 12.767145334803704
      8'hA4: square_root = 8'hCC; // 12.806248474865697
      8'hA5: square_root = 8'hCD; // 12.84523257866513
      8'hA6: square_root = 8'hCE; // 12.884098726725126
      8'hA7: square_root = 8'hCE; // 12.922847983320086
      8'hA8: square_root = 8'hCF; // 12.96148139681572
      8'hA9: square_root = 8'hD0; // 13.0
      8'hAA: square_root = 8'hD0; // 13.038404810405298
      8'hAB: square_root = 8'hD1; // 13.076696830622021
      8'hAC: square_root = 8'hD1; // 13.114877048604
      8'hAD: square_root = 8'hD2; // 13.152946437965905
      8'hAE: square_root = 8'hD3; // 13.19090595827292
      8'hAF: square_root = 8'hD3; // 13.228756555322953
      8'hB0: square_root = 8'hD4; // 13.2664991614216
      8'hB1: square_root = 8'hD4; // 13.30413469565007
      8'hB2: square_root = 8'hD5; // 13.341664064126334
      8'hB3: square_root = 8'hD6; // 13.379088160259652
      8'hB4: square_root = 8'hD6; // 13.416407864998739
      8'hB5: square_root = 8'hD7; // 13.45362404707371
      8'hB6: square_root = 8'hD7; // 13.490737563232042
      8'hB7: square_root = 8'hD8; // 13.527749258468683
      8'hB8: square_root = 8'hD9; // 13.564659966250536
      8'hB9: square_root = 8'hD9; // 13.601470508735444
      8'hBA: square_root = 8'hDA; // 13.638181696985855
      8'hBB: square_root = 8'hDA; // 13.674794331177344
      8'hBC: square_root = 8'hDB; // 13.711309200802088
      8'hBD: square_root = 8'hDB; // 13.74772708486752
      8'hBE: square_root = 8'hDC; // 13.784048752090222
      8'hBF: square_root = 8'hDD; // 13.820274961085254
      8'hC0: square_root = 8'hDD; // 13.856406460551018
      8'hC1: square_root = 8'hDE; // 13.892443989449804
      8'hC2: square_root = 8'hDE; // 13.92838827718412
      8'hC3: square_root = 8'hDF; // 13.96424004376894
      8'hC4: square_root = 8'hE0; // 14.0
      8'hC5: square_root = 8'hE0; // 14.035668847618199
      8'hC6: square_root = 8'hE1; // 14.071247279470288
      8'hC7: square_root = 8'hE1; // 14.106735979665885
      8'hC8: square_root = 8'hE2; // 14.142135623730951
      8'hC9: square_root = 8'hE2; // 14.177446878757825
      8'hCA: square_root = 8'hE3; // 14.212670403551895
      8'hCB: square_root = 8'hE3; // 14.247806848775006
      8'hCC: square_root = 8'hE4; // 14.2828568570857
      8'hCD: square_root = 8'hE5; // 14.317821063276353
      8'hCE: square_root = 8'hE5; // 14.352700094407323
      8'hCF: square_root = 8'hE6; // 14.38749456993816
      8'hD0: square_root = 8'hE6; // 14.422205101855956
      8'hD1: square_root = 8'hE7; // 14.45683229480096
      8'hD2: square_root = 8'hE7; // 14.491376746189438
      8'hD3: square_root = 8'hE8; // 14.52583904633395
      8'hD4: square_root = 8'hE8; // 14.560219778561036
      8'hD5: square_root = 8'hE9; // 14.594519519326424
      8'hD6: square_root = 8'hEA; // 14.628738838327793
      8'hD7: square_root = 8'hEA; // 14.66287829861518
      8'hD8: square_root = 8'hEB; // 14.696938456699069
      8'hD9: square_root = 8'hEB; // 14.730919862656235
      8'hDA: square_root = 8'hEC; // 14.7648230602334
      8'hDB: square_root = 8'hEC; // 14.798648586948742
      8'hDC: square_root = 8'hED; // 14.832396974191326
      8'hDD: square_root = 8'hED; // 14.866068747318506
      8'hDE: square_root = 8'hEE; // 14.89966442575134
      8'hDF: square_root = 8'hEE; // 14.933184523068078
      8'hE0: square_root = 8'hEF; // 14.966629547095765
      8'hE1: square_root = 8'hF0; // 15.0
      8'hE2: square_root = 8'hF0; // 15.033296378372908
      8'hE3: square_root = 8'hF1; // 15.066519173319364
      8'hE4: square_root = 8'hF1; // 15.0996688705415
      8'hE5: square_root = 8'hF2; // 15.132745950421556
      8'hE6: square_root = 8'hF2; // 15.165750888103101
      8'hE7: square_root = 8'hF3; // 15.198684153570664
      8'hE8: square_root = 8'hF3; // 15.231546211727817
      8'hE9: square_root = 8'hF4; // 15.264337522473747
      8'hEA: square_root = 8'hF4; // 15.297058540778355
      8'hEB: square_root = 8'hF5; // 15.329709716755891
      8'hEC: square_root = 8'hF5; // 15.362291495737216
      8'hED: square_root = 8'hF6; // 15.394804318340652
      8'hEE: square_root = 8'hF6; // 15.427248620541512
      8'hEF: square_root = 8'hF7; // 15.459624833740307
      8'hF0: square_root = 8'hF7; // 15.491933384829668
      8'hF1: square_root = 8'hF8; // 15.524174696260024
      8'hF2: square_root = 8'hF8; // 15.556349186104045
      8'hF3: square_root = 8'hF9; // 15.588457268119896
      8'hF4: square_root = 8'hF9; // 15.620499351813308
      8'hF5: square_root = 8'hFA; // 15.652475842498529
      8'hF6: square_root = 8'hFA; // 15.684387141358123
      8'hF7: square_root = 8'hFB; // 15.716233645501712
      8'hF8: square_root = 8'hFB; // 15.748015748023622
      8'hF9: square_root = 8'hFC; // 15.7797338380595
      8'hFA: square_root = 8'hFC; // 15.811388300841896
      8'hFB: square_root = 8'hFD; // 15.84297951775486
      8'hFC: square_root = 8'hFD; // 15.874507866387544
      8'hFD: square_root = 8'hFE; // 15.905973720586866
      8'hFE: square_root = 8'hFE; // 15.937377450509228
      8'hFF: square_root = 8'hFF; // 15.968719422671311
      default: ;
    endcase
  end: ibis_square_root_combinatorial
endmodule: ibis_square_root
